`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    // ROM 크기를 충분히 크게 설정 (256개 엔트리)
    logic [31:0] rom[0:255];

    initial begin
        // R-Type 명령어들 (ALU operations)
        rom[0] = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x2, x1      (12 + 11 = 23)
        rom[1] = 32'b0100000_00001_00010_000_00101_0110011; // sub x5, x2, x1      (12 - 11 = 1)
        rom[2] = 32'b0000000_00001_00010_001_00110_0110011; // sll x6, x2, x1      (12 << 11 = 24576)
        rom[3] = 32'b0000000_00001_00010_010_00111_0110011; // slt x7, x2, x1      (12 < 11 = 0)
        rom[4] = 32'b0000000_00001_00010_011_01000_0110011; // sltu x8, x2, x1     (12 < 11 = 0)
        rom[5] = 32'b0000000_00001_00010_100_01001_0110011; // xor x9, x2, x1      (12 ^ 11 = 7)
        rom[6] = 32'b0000000_00001_00010_101_01010_0110011; // srl x10, x2, x1     (12 >> 11 = 0)
        rom[7] = 32'b0100000_00001_00010_101_01011_0110011; // sra x11, x2, x1     (12 >>> 11 = 0)
        rom[8] = 32'b0000000_00001_00010_110_01100_0110011; // or x12, x2, x1      (12 | 11 = 15)
        rom[9] = 32'b0000000_00001_00010_111_01101_0110011; // and x13, x2, x1     (12 & 11 = 8)

        // I-Type 명령어들 (Immediate ALU operations)
        rom[10] = 32'b000000000101_00010_000_01110_0010011; // addi x14, x2, 5     (12 + 5 = 17)
        rom[11] = 32'b000000100010_00010_010_01111_0010011; // slti x15, x2, 2     (12 < 34 = 1)
        rom[12] = 32'b000000100010_00010_011_10000_0010011; // sltiu x16, x2, 2    (12 < 34 = 1)
        rom[13] = 32'b000000000111_00010_100_10001_0010011; // xori x17, x2, 7     (12 ^ 7 = 11)
        rom[14] = 32'b000000000111_00010_110_10010_0010011; // ori x18, x2, 7      (12 | 7 = 15)
        rom[15] = 32'b000000000111_00010_111_10011_0010011; // andi x19, x2, 7     (12 & 7 = 4)
        rom[16] = 32'b0000000_00010_00010_001_10100_0010011; // slli x20, x2, 2     (12 << 2 = 48)
        rom[17] = 32'b0000000_00010_00010_101_10101_0010011; // srli x21, x2, 2     (12 >> 2 = 3)
        rom[18] = 32'b0100000_00010_00010_101_10110_0010011; // srai x22, x2, 2     (12 >>> 2 = 3)

        // S-Type 명령어들 (Store operations)
        rom[19] = 32'b0000000_00100_00000_010_00100_0100011; // sw x4, 4(x0)        (메모리[4] = x4)
        rom[20] = 32'b0000000_00100_00000_001_01000_0100011; // sh x4, 8(x0)        (메모리[8] = x4의 하위 16비트)
        rom[21] = 32'b0000000_00100_00000_000_01100_0100011; // sb x4, 12(x0)       (메모리[12] = x4의 하위 8비트)

        // L-Type 명령어들 (Load operations)
        rom[22] = 32'b000000000100_00000_010_10111_0000011; // lw x23, 4(x0)       (x23 = 메모리[4] 전체 32비트)
        rom[23] = 32'b000000001000_00000_001_11000_0000011; // lh x24, 8(x0)       (x24 = 메모리[8] 하위 16비트)
        rom[24] = 32'b000000001000_00000_101_11001_0000011; // lhu x25, 8(x0)      (x25 = 메모리[8] 하위 16비트)
        rom[25] = 32'b000000001100_00000_000_11010_0000011; // lb x26, 12(x0)      (x26 = 메모리[12] 하위 8비트)
        rom[26] = 32'b000000001100_00000_100_11011_0000011; // lbu x27, 12(x0)     (x27 = 메모리[12] 하위 8비트)

        // U-Type 명령어들 (Upper immediate) 
        rom[27] = 32'b00000000000000010010_11100_0110111; // lui x28, 0x12        (x28 = 0x12000)
        rom[28] = 32'b00000000000000010010_11101_0010111; // auipc x29, 0x12      (x29 = PC + 0x12000)

        // J-Type 명령어들 (Jump) 
        rom[29] = 32'b0_0000000100_0_00000000_10110_1101111; // jal x22, 4          (x22 = PC+4, PC += 4)
        rom[30] = 32'b000000000000_10110_000_10111_1100111;  // jalr x23, x22, 0    (x23 = PC+4, PC = x22+0)

        for (int i = 31; i < 256; i++) begin
            rom[i] = 32'b000000000000_00000_000_00000_0010011; // addi x0, x0, 0 (NOP)
        end
    end

    assign data = rom[addr[31:2]];
endmodule

